 module test (
  
	input  [4:0] a,b,
	input  [4:0] c,d,
	output  [5:0] result1,
	output  [5:0] result2
);

assign result1=a+b ;
assign result2=c+d ; 

 endmodule 

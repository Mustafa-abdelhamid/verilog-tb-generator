 module test (
	input wire [4:0] a,b,
	output wire [5:0] result
);

assign result=a+b ; 

 endmodule 
